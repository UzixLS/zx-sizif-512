`ifdef REV_C
    `define BANK_PENT_0   4'd0
    `define BANK_S128_0   4'd0
    `define BANK_S128_1   4'd1
    `define BANK_MAGIC    4'd2
    `define BANK_DIV      4'd3
    `define BANK_S3_0     4'd4
    `define BANK_S3_1     4'd5
    `define BANK_S3_2     4'd6
    `define BANK_S3_3     4'd1
    `define BANK_S3_3_DIV 4'd1
    `define BANK_48       4'd1
    `define BANK_48ALT1   4'd7
    `define BANK_48ALT2   4'd7
`else
    `define BANK_PENT_0   4'd0
    `define BANK_S128_0   4'd9
    `define BANK_S128_1   4'd1
    `define BANK_MAGIC    4'd2
    `define BANK_DIV      4'd3
    `define BANK_S3_0     4'd4
    `define BANK_S3_1     4'd5
    `define BANK_S3_2     4'd6
    `define BANK_S3_3     4'd11
    `define BANK_S3_3_DIV 4'd12
    `define BANK_48       4'd10
    `define BANK_48ALT1   4'd7
    `define BANK_48ALT2   4'd8
`endif

import common::*;
module mem(
    input clk28,
    cpu_bus bus,
    inout [7:0] xd,
    output [17:14] ra,
    output reg n_romcs,
    output [18:0] va,
    inout [7:0] vd,
    output n_vrd,
    output reg n_vwr,

    output basic48_paged,

    input machine_t machine,
    input rom_wren,
    input magic_map,
    input [2:0] ram_page128,
    input rom_page128,
    input [2:0] port_1ffd,
    input [4:0] port_dffd,
    input [2:0] ram_pageext,
    input rom_alt48_en,
    input rom_alt48,
    input rom_custom_en,
    input [1:0] rom_custom,
    input divmmc_en,
    input div_ram,
    input div_map,
    input div_ramwr_mask,
    input [3:0] div_page,

    input snow,
    input video_page,
    input video_read_req,
    input video_read_req_is_up,
    input [14:0] video_read_addr,
    input [5:0] video_read_up_addr,
    input up_write_req,
    input [5:0] up_write_addr,

    input magic_dout_active,
    input [7:0] magic_dout,
    input up_dout_active,
    input [7:0] up_dout,
    input div_dout_active,
    input [7:0] div_dout,
    input ay_dout_active,
    input ports_dout_active,
    input [7:0] ports_dout
);

wire [18:13] ram_a;

assign n_vrd = 1'b0;

reg romreq, ramreq;
always @(posedge clk28) begin
    romreq =  bus.mreq && !bus.rfsh && bus.a[15:14] == 2'b00 &&
        (magic_map || (!div_ram && div_map) || (!div_ram && !port_dffd[4] && !port_1ffd[0]));
    ramreq = (bus.mreq && !bus.rfsh && !romreq) || up_write_req;

    n_vwr = ~(ramreq && bus.wr && !div_ramwr_mask && !video_read_req);
    n_romcs = ~romreq;
end

reg vwr0;
reg [7:0] xd_bufwr;
reg [18:0] va_buf;
always @(negedge clk28) begin
    if (~n_vwr && !vwr0)
        xd_bufwr <= xd;
    vwr0 <= ~n_vwr;

    if (bus.mreq && ramreq)
        va_buf <= {ram_a[18:13], bus.a[12:0]};
end


// reserve 128K RAM for DivMMC
wire [1:0] ram_pageext0 = {divmmc_en? 1'b1 : ~ram_pageext[1], ~ram_pageext[0]};

assign ram_a =
    (magic_map && bus.a[15:14] == 2'b11)           ? {2'b00, 3'b111, bus.a[13]} :
    (magic_map)                                    ? {3'b111, video_page, bus.a[14:13]} :
    (div_map && bus.a[15:13] == 3'b001)            ? {2'b01, div_page} :
    (div_map && bus.a[15:14] == 2'b00)             ? {2'b01, 4'b0011} :
    (port_dffd[3] && bus.a[15])                    ? {2'b11, bus.a[14], bus.a[15], bus.a[14], bus.a[13]} :
    (port_dffd[3] && bus.a[14])                    ? {ram_pageext0, ram_page128, bus.a[13]} :
    (port_1ffd[2] == 1'b0 && port_1ffd[0] == 1'b1) ? {2'b11, port_1ffd[1], bus.a[15], bus.a[14], bus.a[13]} :
    (port_1ffd == 3'b101)                          ? {2'b11, ~(bus.a[15] & bus.a[14]), bus.a[15], bus.a[14], bus.a[13]} :
    (port_1ffd == 3'b111)                          ? {2'b11, ~(bus.a[15] & bus.a[14]), (bus.a[15] | bus.a[14]), bus.a[14], bus.a[13]} :
    (bus.a[15:14] == 2'b11)                        ? {ram_pageext0, ram_page128, bus.a[13]} :
                                                     {2'b11, bus.a[14], bus.a[15], bus.a[14], bus.a[13]} ;


assign ra[17:14] =
    rom_wren                                          ? {3'b000, bus.a[0]} : // handle jedec sequence (Z80 addr #1555 = ROM addr #05555, Z80 addr #2AAA = ROM addr #02AAA)
    magic_map                                         ? `BANK_MAGIC :
    div_map                                           ? `BANK_DIV :
`ifndef REV_C
    (rom_custom_en && rom_page128 == 1'b0)            ? {2'b11, rom_custom} :
`endif
    (machine == MACHINE_S3)? (
        (port_1ffd[2] == 1'b0 && rom_page128 == 1'b0) ? `BANK_S3_0 :
        (port_1ffd[2] == 1'b0 && rom_page128 == 1'b1) ? `BANK_S3_1 :
        (port_1ffd[2] == 1'b1 && rom_page128 == 1'b0) ? `BANK_S3_2 :
        (rom_alt48_en && rom_alt48)                   ? `BANK_48ALT2 :
        (rom_alt48_en)                                ? `BANK_48ALT1 :
        (divmmc_en)                                   ? `BANK_S3_3_DIV :
                                                        `BANK_S3_3 ) :
    (machine == MACHINE_S128)? (
        (rom_page128 == 1'b0)                         ? `BANK_S128_0 :
        (rom_alt48_en && rom_alt48)                   ? `BANK_48ALT2 :
        (rom_alt48_en)                                ? `BANK_48ALT1 :
                                                        `BANK_S128_1 ) :
    (machine == MACHINE_PENT)? (
        (rom_page128 == 1'b0)                         ? `BANK_PENT_0 :
        (rom_alt48_en && rom_alt48)                   ? `BANK_48ALT2 :
        (rom_alt48_en)                                ? `BANK_48ALT1 :
                                                        `BANK_S128_1 ) :
    // 48K
    (rom_alt48_en && rom_alt48)                       ? `BANK_48ALT2 :
    (rom_alt48_en)                                    ? `BANK_48ALT1 :
                                                        `BANK_48 ;

assign basic48_paged = (ra == `BANK_48) ||
                       (ra == `BANK_48ALT1) ||
                       (ra == `BANK_48ALT2) ||
                       (ra == `BANK_S128_1) ||
                       (ra == `BANK_S3_3) ||
                       (ra == `BANK_S3_3_DIV) ;


assign va[18:0] =
    video_read_req && video_read_req_is_up ? {2'b00, 3'b111, 8'b11111111, video_read_up_addr} :
    video_read_req && snow                 ? {3'b111, video_page, video_read_addr[14:8], bus.a[7:0]} :
    video_read_req                         ? {3'b111, video_page, video_read_addr} :
    up_write_req                           ? {2'b00, 3'b111, 8'b11111111, up_write_addr} :
                                             va_buf;


// this is required because of weak xd pullup causing garbage reads from nonexisting ports
reg [1:0] xd_precharge0;
wire xd_precharge = clk28 && xd_precharge0[1] && !xd_precharge0[0];
always @(posedge clk28)
    xd_precharge0 <= {bus.iorq && (bus.rd || bus.m1), xd_precharge0[1]};

assign xd[7:0] =
    (ramreq && bus.rd)             ? vd :
    magic_dout_active              ? magic_dout :
    up_dout_active                 ? up_dout :
    div_dout_active                ? div_dout :
    ay_dout_active                 ? {8{1'bz}} :
    ports_dout_active              ? ports_dout :
    xd_precharge                   ? 8'hFF :
                                     {8{1'bz}} ;

assign vd[7:0] =
    (~n_vwr & vwr0)                ? xd_bufwr :
                                     {8{1'bz}} ;


endmodule
