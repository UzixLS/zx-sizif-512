// A-Z
`define PS2_A           9'h1C
`define PS2_B           9'h32
`define PS2_C           9'h21
`define PS2_D           9'h23
`define PS2_E           9'h24
`define PS2_F           9'h2B
`define PS2_G           9'h34
`define PS2_H           9'h33
`define PS2_I           9'h43
`define PS2_J           9'h3B
`define PS2_K           9'h42
`define PS2_L           9'h4B
`define PS2_M           9'h3A
`define PS2_N           9'h31
`define PS2_O           9'h44
`define PS2_P           9'h4D
`define PS2_Q           9'h15
`define PS2_R           9'h2D
`define PS2_S           9'h1B
`define PS2_T           9'h2C
`define PS2_U           9'h3C
`define PS2_V           9'h2A
`define PS2_W           9'h1D
`define PS2_X           9'h22
`define PS2_Y           9'h35
`define PS2_Z           9'h1A

// 0-9
`define PS2_0           9'h45
`define PS2_1           9'h16
`define PS2_2           9'h1E
`define PS2_3           9'h26
`define PS2_4           9'h25
`define PS2_5           9'h2E
`define PS2_6           9'h36
`define PS2_7           9'h3D
`define PS2_8           9'h3E
`define PS2_9           9'h46

// Others
`define PS2_ACCENT      9'h0E    // '`'
`define PS2_MINUS       9'h4E    // '-'
`define PS2_EQUALS      9'h55    // '='
`define PS2_BACK_SLASH  9'h5D    // '\'
`define PS2_SPACE       9'h29    // ' '
`define PS2_TAB         9'h0D    // '\t'
`define PS2_L_BRACKET   9'h54    // '['
`define PS2_R_BRACKET   9'h5B    // ']'
`define PS2_SEMICOLON   9'h4C    // ';'
`define PS2_QUOTE       9'h52    // '''
`define PS2_COMMA       9'h41    // ','
`define PS2_PERIOD      9'h49    // '.'
`define PS2_SLASH       9'h4A    // '/'

// Control
`define PS2_BACKSPACE   9'h66
`define PS2_CAPS        9'h58
`define PS2_SCROLL      9'h7E
`define PS2_NUM         9'h77
`define PS2_L_SHIFT     9'h12
`define PS2_R_SHIFT     9'h59
`define PS2_L_CTRL      9'h14
`define PS2_R_CTRL      9'h114
`define PS2_L_ALT       9'h11
`define PS2_R_ALT       9'h111
`define PS2_ENTER       9'h5A
`define PS2_ESC         9'h76
`define PS2_INSERT      9'h170
`define PS2_DELETE      9'h171
`define PS2_HOME        9'h16C
`define PS2_END         9'h169
`define PS2_PGUP        9'h17D
`define PS2_PGDN        9'h17A
`define PS2_UP          9'h175
`define PS2_DOWN        9'h172
`define PS2_LEFT        9'h16B
`define PS2_RIGHT       9'h174
`define PS2_PSCR1       9'h112
`define PS2_PSCR2       9'h17c
`define PS2_L_WIN       9'h11f
`define PS2_R_WIN       9'h127
`define PS2_MENU        9'h12f
`define PS2_PAUSE       9'h177


// F1..F12
`define PS2_F1          9'h05
`define PS2_F2          9'h06
`define PS2_F3          9'h04
`define PS2_F4          9'h0C
`define PS2_F5          9'h03
`define PS2_F6          9'h0B
`define PS2_F7          9'h83
`define PS2_F8          9'h0A
`define PS2_F9          9'h01
`define PS2_F10         9'h09
`define PS2_F11         9'h78
`define PS2_F12         9'h07

// Keypad
`define PS2_NUMLOCK     9'h77
`define PS2_KP_SLASH    9'h14A
`define PS2_KP_STAR     9'h7C
`define PS2_KP_MINUS    9'h7B
`define PS2_KP_PLUS     9'h79
`define PS2_KP_ENTER    9'h15A
`define PS2_KP_PERIOD   9'h71
`define PS2_KP_0        9'h70
`define PS2_KP_1        9'h69
`define PS2_KP_2        9'h72
`define PS2_KP_3        9'h7A
`define PS2_KP_4        9'h6B
`define PS2_KP_5        9'h73
`define PS2_KP_6        9'h74
`define PS2_KP_7        9'h6C
`define PS2_KP_8        9'h75
`define PS2_KP_9        9'h7D

